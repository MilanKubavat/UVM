package ClockResetPkg;

  `include "uvm_macros.svh"

  import uvm_pkg::*;

  `include "ClockResetCfg.sv"

  `include "ClockDriver.sv"
  `include "ClockMonitor.sv"
  `include "ClockAgent.sv"

  `include "ResetDriver.sv"
  `include "ResetMonitor.sv"
  `include "ResetAgent.sv"

  `include "ClockResetEnv.sv"

  `include "ClockResetBaseTest.sv"

endpackage
