//----------------------------------------------------------
// Start Date: 10 Apr 2020
// Last Modified:
// Author: Milan Kubavat
// 
// Description: ahb master pkg to compile ahb master 
//----------------------------------------------------------

package ahb_master_pkg;

  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import ahb_common_pkg::*;

  `include "ahb_master_cfg.sv"
  `include "ahb_master_seq_lib.sv"
  `include "ahb_master_sequencer.sv"
  `include "ahb_master_driver.sv"
  `include "ahb_master_agent.sv"

endpackage
