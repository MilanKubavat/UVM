//----------------------------------------------------------
// Start Date: 10 Apr 2020
// Last Modified:
// Author: Milan Kubavat
// 
// Description: AMBA3 AHB-Lite interface
//----------------------------------------------------------

interface ahb_interface (input HCLK, HRESETn);
endinterface	
